module main

// Stub methods for parser submodules.
// All declaration stubs have been moved to declarations.v.
// This file is kept for any remaining stubs from untranslated files.
